* File: inv.pex.netlist
* Created: Tue Nov  4 23:53:44 2025
* Program "Calibre xRC"
* Version "v2024.4_12.9"
* 
.include "inv.pex.netlist.pex"
.subckt inv  GND! OUT VDD! A1
* 
* A1	A1
* VDD!	VDD!
* INV	INV
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=5.12015e-12
+ PERIM=9.142e-06
XMMN0 N_OUT_MMN0_d N_A1_MMN0_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET L=6.8e-08
+ W=1e-06 AD=5.51e-13 AS=5.51e-13 PD=3.102e-06 PS=3.102e-06 NRD=0.382 NRS=0.382
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=5.51e-07 SB=5.51e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=4.692e-15 PANW8=1.36e-14
+ PANW9=2.72e-14 PANW10=2.2508e-14
XMMP0 N_OUT_MMP0_d N_A1_MMP0_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET L=6.8e-08
+ W=1.3e-06 AD=7.163e-13 AS=7.163e-13 PD=3.702e-06 PS=3.702e-06 NRD=0.293846
+ NRS=0.293846 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=5.51e-07
+ SB=5.51e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.264e-15 PANW6=6.8e-15
+ PANW7=1.36e-14 PANW8=1.1186e-13 PANW9=1.428e-13 PANW10=6.4736e-14
*
.include "inv.pex.netlist.INV.pxi"
*
.ends
*
*
